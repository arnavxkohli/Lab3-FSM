module clktick #(
)(
  // interface signals
);

endmodule
